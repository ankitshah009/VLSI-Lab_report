magic
tech scmos
timestamp 1395901728
<< nwell >>
rect -4 16 17 27
<< polysilicon >>
rect 1 27 3 29
rect 10 27 12 29
rect 1 -1 3 16
rect 10 -1 12 16
rect 1 -7 3 -5
rect 10 -7 12 -5
<< ndiffusion >>
rect 0 -5 1 -1
rect 3 -5 10 -1
rect 12 -5 13 -1
<< pdiffusion >>
rect 0 23 1 27
rect -4 16 1 23
rect 3 20 10 27
rect 3 16 4 20
rect 8 16 10 20
rect 12 23 13 27
rect 12 16 17 23
<< metal1 >>
rect -4 33 17 42
rect -4 27 0 33
rect 13 27 17 33
rect 4 5 8 16
rect 4 1 17 5
rect 13 -1 17 1
rect -4 -11 0 -5
rect -4 -19 18 -11
<< ntransistor >>
rect 1 -5 3 -1
rect 10 -5 12 -1
<< ptransistor >>
rect 1 16 3 27
rect 10 16 12 27
<< polycontact >>
rect -3 8 1 12
rect 12 9 16 13
<< ndcontact >>
rect -4 -5 0 -1
rect 13 -5 17 -1
<< pdcontact >>
rect -4 23 0 27
rect 4 16 8 20
rect 13 23 17 27
<< labels >>
rlabel metal1 5 37 5 37 5 vdd
<< end >>
