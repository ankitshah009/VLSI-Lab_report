magic
tech scmos
timestamp 1397105118
<< nwell >>
rect -18 14 13 42
<< polysilicon >>
rect -12 25 -10 27
rect -3 25 -1 27
rect 6 25 8 27
rect -12 -3 -10 15
rect -3 -3 -1 15
rect 6 -3 8 15
rect -12 -9 -10 -7
rect -3 -9 -1 -7
rect 6 -9 8 -7
<< ndiffusion >>
rect -13 -7 -12 -3
rect -10 -7 -8 -3
rect -4 -7 -3 -3
rect -1 -7 0 -3
rect 4 -7 6 -3
rect 8 -7 9 -3
<< pdiffusion >>
rect -13 22 -12 25
rect -17 19 -12 22
rect -13 15 -12 19
rect -10 21 -8 25
rect -4 21 -3 25
rect -10 18 -3 21
rect -10 15 -8 18
rect -4 15 -3 18
rect -1 15 6 25
rect 8 22 9 25
rect 8 19 13 22
rect 8 15 9 19
<< metal1 >>
rect -8 38 9 42
rect -8 34 13 38
rect -17 19 -13 22
rect -17 -3 -13 15
rect -8 25 -4 34
rect -8 18 -4 21
rect 9 19 13 22
rect 9 6 13 15
rect 0 4 13 6
rect -6 3 13 4
rect -6 0 4 3
rect 0 -3 4 0
rect -8 -12 -4 -7
rect 9 -12 13 -7
rect -8 -19 13 -12
<< ntransistor >>
rect -12 -7 -10 -3
rect -3 -7 -1 -3
rect 6 -7 8 -3
<< ptransistor >>
rect -12 15 -10 25
rect -3 15 -1 25
rect 6 15 8 25
<< polycontact >>
rect -7 7 -3 11
rect -10 0 -6 4
rect 2 9 6 13
<< ndcontact >>
rect -17 -7 -13 -3
rect -8 -7 -4 -3
rect 0 -7 4 -3
rect 9 -7 13 -3
<< pdcontact >>
rect -17 22 -13 26
rect -17 15 -13 19
rect -8 21 -4 25
rect -8 14 -4 18
rect 9 22 13 26
rect 9 15 13 19
<< nsubstratencontact >>
rect 9 38 13 42
<< labels >>
rlabel metal1 2 -15 2 -15 1 vss
rlabel metal1 1 38 1 38 5 vdd
rlabel polycontact 4 11 4 11 1 b
rlabel pdiffusion 3 21 3 21 1 d1s2p
rlabel polycontact -5 9 -5 9 1 a
rlabel metal1 -15 6 -15 6 3 out
rlabel metal1 11 8 11 8 7 out1
<< end >>
