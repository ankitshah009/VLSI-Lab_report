magic
tech scmos
timestamp 1395292474
<< polysilicon >>
rect 11 19 17 21
rect 11 2 17 14
rect 11 -5 17 -3
<< ndiffusion >>
rect 10 -3 11 2
rect 17 -3 18 2
<< pdiffusion >>
rect 10 14 11 19
rect 17 14 18 19
<< metal1 >>
rect 6 22 21 26
rect 6 19 10 22
rect 18 2 22 14
<< metal2 >>
rect 6 -6 10 2
rect 6 -10 21 -6
<< ntransistor >>
rect 11 -3 17 2
<< ptransistor >>
rect 11 14 17 19
<< polycontact >>
rect 6 7 11 11
<< ndcontact >>
rect 6 -3 10 2
rect 18 -3 22 2
<< pdcontact >>
rect 6 14 10 19
rect 18 14 22 19
<< end >>
