

.include /home/krunal/VLSI_LAB/VINAY/t14y_tsmc_025_level3.txt
m1 drn gate s 0 cmosn l=1u w=.5u

vdd drn 0 5
vin gate 0 5
vss s 0 0

.dc  vin 0 6 .1 vss 0 3 1
.control
run 
plot -vdd#branch
.end
