magic
tech scmos
timestamp 1398186171
<< nwell >>
rect -4 16 17 37
<< polysilicon >>
rect 1 27 3 29
rect 10 27 12 29
rect 1 -1 3 16
rect 10 -1 12 16
rect 1 -7 3 -5
rect 10 -7 12 -5
<< ndiffusion >>
rect 0 -5 1 -1
rect 3 -5 10 -1
rect 12 -5 13 -1
<< pdiffusion >>
rect 0 16 1 27
rect 3 20 10 27
rect 3 16 4 20
rect 8 16 10 20
rect 12 16 13 27
<< metal1 >>
rect -4 37 17 42
rect -4 33 13 37
rect -4 27 0 33
rect 13 27 17 33
rect 4 5 8 16
rect 4 1 17 5
rect 13 -1 17 1
rect -4 -11 0 -5
rect -4 -19 18 -11
<< ntransistor >>
rect 1 -5 3 -1
rect 10 -5 12 -1
<< ptransistor >>
rect 1 16 3 27
rect 10 16 12 27
<< polycontact >>
rect -3 8 1 12
rect 12 9 16 13
<< ndcontact >>
rect -4 -5 0 -1
rect 13 -5 17 -1
<< pdcontact >>
rect -4 16 0 27
rect 4 16 8 20
rect 13 16 17 27
<< nsubstratencontact >>
rect 13 33 17 37
<< labels >>
rlabel metal1 15 3 15 3 7 out
rlabel polycontact -1 10 -1 10 3 a
rlabel polycontact 14 11 14 11 7 b
rlabel metal1 7 -15 7 -15 1 vss
rlabel ntransistor 2 -3 2 -3 1 nmos1
rlabel ntransistor 11 -3 11 -3 1 nmos2
rlabel ndiffusion 7 -3 7 -3 1 s2d1n
rlabel pdiffusion 6 24 6 24 1 d1d2p
rlabel ptransistor 11 21 11 21 1 pmos2
rlabel ptransistor 2 22 2 22 1 pmos1
rlabel metal1 5 37 5 37 5 vdd
<< end >>
