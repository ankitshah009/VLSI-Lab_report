magic
tech scmos
timestamp 1396498188
<< nwell >>
rect 4 13 19 27
<< polysilicon >>
rect 11 19 13 21
rect 11 2 13 14
rect 11 -5 13 -3
<< ndiffusion >>
rect 10 -3 11 2
rect 13 -3 14 2
<< pdiffusion >>
rect 10 14 11 19
rect 13 14 14 19
<< metal1 >>
rect 6 23 14 26
rect 6 22 18 23
rect 6 19 10 22
rect 14 2 18 14
rect 6 -6 10 -3
rect 6 -10 18 -6
<< ntransistor >>
rect 11 -3 13 2
<< ptransistor >>
rect 11 14 13 19
<< polycontact >>
rect 6 7 11 11
<< ndcontact >>
rect 6 -3 10 2
rect 14 -3 18 2
<< pdcontact >>
rect 6 14 10 19
rect 14 14 18 19
<< nsubstratencontact >>
rect 14 23 18 27
<< labels >>
rlabel polycontact 8 9 8 9 3 input
rlabel metal1 14 -7 14 -7 1 vss
rlabel metal1 16 8 16 8 7 out
rlabel metal1 14 24 14 24 5 vdd
<< end >>
