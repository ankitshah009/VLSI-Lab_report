magic
tech scmos
timestamp 1398193493
<< nwell >>
rect -8 14 13 38
<< polysilicon >>
rect -3 25 -1 27
rect 6 25 8 27
rect -3 -3 -1 15
rect 6 -3 8 15
rect -3 -9 -1 -7
rect 6 -9 8 -7
<< ndiffusion >>
rect -4 -7 -3 -3
rect -1 -7 0 -3
rect 4 -7 6 -3
rect 8 -7 9 -3
<< pdiffusion >>
rect -4 15 -3 25
rect -1 15 6 25
rect 8 15 9 25
<< metal1 >>
rect -8 34 9 38
rect -8 30 13 34
rect -8 25 -4 30
rect 9 6 13 15
rect 0 3 13 6
rect 0 -3 4 3
rect -8 -12 -4 -7
rect 9 -12 13 -7
rect -8 -19 13 -12
<< ntransistor >>
rect -3 -7 -1 -3
rect 6 -7 8 -3
<< ptransistor >>
rect -3 15 -1 25
rect 6 15 8 25
<< polycontact >>
rect -7 7 -3 11
rect 2 9 6 13
<< ndcontact >>
rect -8 -7 -4 -3
rect 0 -7 4 -3
rect 9 -7 13 -3
<< pdcontact >>
rect -8 15 -4 25
rect 9 15 13 26
<< nsubstratencontact >>
rect 9 34 13 38
<< labels >>
rlabel metal1 2 -15 2 -15 1 vss
rlabel polycontact 4 11 4 11 1 b
rlabel pdiffusion 3 21 3 21 1 d1s2p
rlabel polycontact -5 9 -5 9 1 a
rlabel metal1 11 8 11 8 7 out1
rlabel metal1 1 34 1 34 5 vdd
<< end >>
